// Modified by Princeton University on June 9th, 2015
// ========== Copyright Header Begin ==========================================
//
// OpenSPARC T1 Processor File: cmp_top.v
// Copyright (c) 2006 Sun Microsystems, Inc.  All Rights Reserved.
// DO NOT ALTER OR REMOVE COPYRIGHT NOTICES.
//
// The above named program is free software; you can redistribute it and/or
// modify it under the terms of the GNU General Public
// License version 2 as published by the Free Software Foundation.
//
// The above named program is distributed in the hope that it will be
// useful, but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
// General Public License for more details.
//
// You should have received a copy of the GNU General Public
// License along with this work; if not, write to the Free Software
// Foundation, Inc., 51 Franklin St, Fifth Floor, Boston, MA 02110-1301, USA.
//
// ========== Copyright Header End ============================================
////////////////////////////////////////////////////////

`ifndef USE_TEST_TOP // don't compile if user wants to use deprecated TOPs
`include "sys.h"
`include "iop.h"
`include "cross_module.tmp.h"
`include "ifu.tmp.h"
`include "define.tmp.h"
`include "piton_system.vh"
`include "jtag.vh"


// /home/alireza/work/git/OpenPiton/OpenPiton-Mess-integration/piton/verif/env/manycore/devices_ariane.xml




`ifdef PITON_DPI
import "DPI-C" function longint read_64b_call (input longint addr);
import "DPI-C" function void write_64b_call (input longint addr, input longint data);
import "DPI-C" function int drive_iob ();
import "DPI-C" function int get_cpx_word (int index);
import "DPI-C" function void report_pc (longint thread_pc);
import "DPI-C" function void init_jbus_model_call(string str, int oram);

`ifndef VERILATOR
// MPI Yummy functions
import "DPI-C" function void initialize();
import "DPI-C" function void finalize();
import "DPI-C" function int getRank();
import "DPI-C" function int getSize();

import "DPI-C" function void mpi_send_yummy(input byte unsigned message, input int dest, input int rank, input int flag);
import "DPI-C" function byte unsigned mpi_receive_yummy(input int origin, input int flag);

import "DPI-C" function longint unsigned mpi_receive_data(input int origin, output byte unsigned valid, input int flag);
import "DPI-C" function void mpi_send_data(input longint unsigned data, input byte unsigned valid, input int dest, input int rank, input int flag);

import "DPI-C" function void barrier();
//add metro_stuff
`endif // ifndef VERILATOR
`endif // ifdef PITON_DPI






`timescale 1ps/1ps
module metro_chipset (
`ifdef VERILATOR
	core_ref_clk,

	sys_rst_n,

	pll_rst_n,

	clk_en,

	pll_bypass,
	pll_rangea,
	pll_lock,
	clk_mux_sel,
	async_mux,
	diag_done,
	ok_iob,

	noc_chanel_in	,
	noc_chanel_out	,
	smart_max,
    flit_o_cnts,
    flit_i_cnts,

/*
input wire                            processor_offchip_noc1_valid,
input wire [`NOC_DATA_WIDTH-1:0]    processor_offchip_noc1_data,
output wire                           processor_offchip_noc1_yummy,
input wire                            processor_offchip_noc2_valid,
input wire [`NOC_DATA_WIDTH-1:0]    processor_offchip_noc2_data,
output wire                           processor_offchip_noc2_yummy,
input wire                            processor_offchip_noc3_valid,
input wire [`NOC_DATA_WIDTH-1:0]    processor_offchip_noc3_data,
output wire                           processor_offchip_noc3_yummy,

output wire                           offchip_processor_noc1_valid,
output wire [`NOC_DATA_WIDTH-1:0]   offchip_processor_noc1_data,
input  wire                           offchip_processor_noc1_yummy,
output wire                           offchip_processor_noc2_valid,
output wire [`NOC_DATA_WIDTH-1:0]   offchip_processor_noc2_data,
input  wire                           offchip_processor_noc2_yummy,
output wire                           offchip_processor_noc3_valid,
output wire [`NOC_DATA_WIDTH-1:0]   offchip_processor_noc3_data,
input  wire                           offchip_processor_noc3_yummy,
*/

	good_end,
	bad_end,
	test_ena
`endif
);


`ifdef PITON_PRONOC
	`include "pronoc_def.v"
 	`NOC_CONF
	
	typedef struct packed {	
		smartflit_chanel_t  [2:0] smartflit_chanel;  		
	} noc_chanel_t;

`else

	typedef struct packed {	
		logic  [`NOC_DATA_WIDTH-1:0] data1;
		logic  [`NOC_DATA_WIDTH-1:0] data2;
		logic  [`NOC_DATA_WIDTH-1:0] data3;
		logic  [2:0] valid;
		logic  [2:0] yummy;		
	} noc_chanel_t;

`endif

localparam NOC_CHANEL_w = $bits(noc_chanel_t); 	


`ifdef VERILATOR

input reg                             core_ref_clk;
input reg                             sys_rst_n;
input reg                             pll_rst_n;
input reg                             clk_en;
input reg                             pll_bypass;
input reg [4:0]                       pll_rangea;
output wire                           pll_lock;
input reg [1:0]                       clk_mux_sel;
input reg                             async_mux;
input                                 diag_done;
input                                 ok_iob;

input  noc_chanel_t noc_chanel_in;
output noc_chanel_t noc_chanel_out;
output [31 : 0] smart_max;
output [63 : 0]   flit_o_cnts,flit_i_cnts;


output wire                           good_end;
output wire                           bad_end;
input  wire                           test_ena;
`endif









//////////////////////
// Type Declarations
//////////////////////

`ifndef VERILATOR
reg                             core_ref_clk;
reg                             sys_rst_n;
reg                             pll_rst_n;
reg                             clk_en;
reg                             pll_bypass;
reg [4:0]                       pll_rangea;
wire                            pll_lock = 1'b1;
reg [1:0]                       clk_mux_sel;
reg                             async_mux;
// For simulation only, monitor stuff.  Only cross-module referenced
// do not delete.
reg                             diag_done;
`endif // ifndef VERILATOR

reg                             io_clk;
reg                             jtag_clk;
reg                             chipset_clk_osc_p;
reg                             chipset_clk_osc_n;
reg                             chipset_clk_osc;
reg                             chipset_clk;
reg                             mem_clk;
reg                             spi_sys_clk;
reg                             chipset_passthru_clk_p;
reg                             chipset_passthru_clk_n;
reg                             passthru_clk_osc_p;
reg                             passthru_clk_osc_n;
reg                             passthru_chipset_clk_p;
reg                             passthru_chipset_clk_n;

reg                             jtag_rst_l;

reg                             jtag_modesel;
reg                             jtag_datain;
wire                            jtag_dataout;


// For simulation only, monitor stuff.  Only cross-module referenced
// do not delete.
reg                             fail_flag;
reg [3:0]                       stub_done;
reg [3:0]                       stub_pass;

`ifndef VERILATOR
reg                       processor_offchip_noc1_valid;
reg [`NOC_DATA_WIDTH-1:0] processor_offchip_noc1_data;
reg                       processor_offchip_noc1_yummy;
reg                       processor_offchip_noc2_valid;
reg [`NOC_DATA_WIDTH-1:0] processor_offchip_noc2_data;
reg                       processor_offchip_noc2_yummy;
reg                       processor_offchip_noc3_valid;
reg [`NOC_DATA_WIDTH-1:0] processor_offchip_noc3_data;
reg                       processor_offchip_noc3_yummy;

reg                       offchip_processor_noc1_valid;
reg [`NOC_DATA_WIDTH-1:0] offchip_processor_noc1_data;
reg                       offchip_processor_noc1_yummy;
reg                       offchip_processor_noc2_valid;
reg [`NOC_DATA_WIDTH-1:0] offchip_processor_noc2_data;
reg                       offchip_processor_noc2_yummy;
reg                       offchip_processor_noc3_valid;
reg [`NOC_DATA_WIDTH-1:0] offchip_processor_noc3_data;
reg                       offchip_processor_noc3_yummy;

`else 

wire                            processor_offchip_noc1_valid;
wire [`NOC_DATA_WIDTH-1:0]      processor_offchip_noc1_data;
wire                            processor_offchip_noc1_yummy;
wire                            processor_offchip_noc2_valid;
wire [`NOC_DATA_WIDTH-1:0]      processor_offchip_noc2_data;
wire                            processor_offchip_noc2_yummy;
wire                            processor_offchip_noc3_valid;
wire [`NOC_DATA_WIDTH-1:0]      processor_offchip_noc3_data;
wire                            processor_offchip_noc3_yummy;

wire                            offchip_processor_noc1_valid;
wire [`NOC_DATA_WIDTH-1:0]      offchip_processor_noc1_data;
wire                            offchip_processor_noc1_yummy;
wire                            offchip_processor_noc2_valid;
wire [`NOC_DATA_WIDTH-1:0]      offchip_processor_noc2_data;
wire                            offchip_processor_noc2_yummy;
wire                            offchip_processor_noc3_valid;
wire [`NOC_DATA_WIDTH-1:0]      offchip_processor_noc3_data;
wire                            offchip_processor_noc3_yummy;



`endif // VERILATOR

////////////////////
// Simulated Clocks
////////////////////

`ifndef VERILATOR
`ifndef USE_FAKE_PLL_AND_CLKMUX
always #5000 core_ref_clk = ~core_ref_clk;                      // 100MHz
`else
always #500 core_ref_clk = ~core_ref_clk;                       // 1000MHz
`endif
`endif

`ifndef VERILATOR
`ifndef SYNC_MUX
always #1429 io_clk = ~io_clk;                                  // 350MHz
`else
always @ * io_clk = core_ref_clk;
`endif
`endif

`ifndef VERILATOR
always #50000 jtag_clk = ~jtag_clk;                             // 10MHz

always #2500 chipset_clk_osc_p = ~chipset_clk_osc_p;            // 200MHz
always @ * chipset_clk_osc_n = ~chipset_clk_osc_p;

always #5000 chipset_clk_osc = ~chipset_clk_osc;                // 100MHz

always #2500 chipset_clk = ~chipset_clk;                        // 200MHz

always #3333 passthru_clk_osc_p = ~passthru_clk_osc_p;          // 150MHz
always @ * passthru_clk_osc_n = ~passthru_clk_osc_p;

always #1429 passthru_chipset_clk_p = ~passthru_chipset_clk_p;  // 350MHz
always @ * passthru_chipset_clk_n = ~passthru_chipset_clk_p;

always #1000 mem_clk = ~mem_clk;                                // 500MHz

always #25000 spi_sys_clk = ~spi_sys_clk;                       // 20MHz
`else

always @(*)    chipset_clk = core_ref_clk;

`endif


initial begin 
 $display("Cache Configuration:");
 $display("\tL2   size:%d,\t associativity:%d",`L2_SIZE,`L2_WAYS);
 $display("\tL1.5 size:%d,\t associativity:%d",`CONFIG_L15_SIZE,`CONFIG_L15_ASSOCIATIVITY);
 $display("\tL1D  size:%d,\t associativity:%d",`CONFIG_L1D_SIZE,`CONFIG_L1D_ASSOCIATIVITY);
 $display("\tL1I  size:%d,\t associativity:%d",`CONFIG_L1I_SIZE,`CONFIG_L1I_ASSOCIATIVITY);
 
 $display("NoC Configuration:");
 $display("\tNOC1 Width:%d",`NOC_DATA_WIDTH);
 $display("\tNOC2 Width:%d",`NOC_DATA_WIDTH);
 $display("\tNOC3 Width:%d",`NOC_DATA_WIDTH);
`ifdef PITON_NO_CHIP_BRIDGE
    $display("**Warning: Chip Bridge Disable"); 
    $display("\t     Only one clock is used in the system"); 
    $display("Clock frequency = 1000 MHz"); 
`endif // PITON_NO_CHIP_BRIDGE
end



////////////////////////////////////////////////////////
// SIMULATED BOOT SEQUENCE
////////////////////////////////////////////////////////

int rank;
int size;
int dest;
byte unsigned valid_aux;

int YUMMY_NOC_1 ;
int DATA_NOC_1  ;
int YUMMY_NOC_2 ;
int DATA_NOC_2  ;
int YUMMY_NOC_3 ;
int DATA_NOC_3  ;

`ifndef VERILATOR
initial
begin
    $dumpfile("metro_chipset.vcd");
    $dumpvars(0, metro_chipset);

    YUMMY_NOC_1 = 0;
    DATA_NOC_1  = 1;
    YUMMY_NOC_2 = 2;
    DATA_NOC_2  = 3;
    YUMMY_NOC_3 = 4;
    DATA_NOC_3  = 5;

    //metro initialization
    initialize();
    //barrier();
    rank = getRank();
    size = getSize();
    $display("METRO_CHIPSET INITIALIZING...");
    $display("size: %d", size);
    $display("rank: %d", rank);
    if (rank==0) begin
            dest = 1;
    end else begin
            dest = 0;
    end
    // These are not referenced elsewhere in this module,
    // but are cross referenced from monitor.v.pyv.  Do not
    // delete
    fail_flag = 1'b0;
    stub_done = 4'b0;
    stub_pass = 4'b0;

    // Clocks initial value
    core_ref_clk = 1'b0;
    io_clk = 1'b0;
    jtag_clk = 1'b0;
    chipset_clk_osc_p = 1'b0;
    chipset_clk_osc_n = 1'b1;
    chipset_clk_osc = 1'b0;
    chipset_clk = 1'b0;
    mem_clk = 1'b0;
    spi_sys_clk = 1'b0;
    chipset_passthru_clk_p = 1'b0;
    chipset_passthru_clk_n = 1'b1;
    passthru_clk_osc_p = 1'b0;
    passthru_clk_osc_n = 1'b1;
    passthru_chipset_clk_p = 1'b0;
    passthru_chipset_clk_n = 1'b1;

    // Resets are held low at start of boot
    sys_rst_n = 1'b0;
    jtag_rst_l = 1'b0;
    pll_rst_n = 1'b0;

    // Mostly DC signals set at start of boot
    clk_en = 1'b0;
    if ($test$plusargs("pll_en"))
    begin
        // PLL is disabled by default
        pll_bypass = 1'b0; // trin: pll_bypass is a switch in the pll; not reliable
        clk_mux_sel[1:0] = 2'b10; // selecting pll
    end
    else
    begin
        pll_bypass = 1'b1; // trin: pll_bypass is a switch in the pll; not reliable
        clk_mux_sel[1:0] = 2'b00; // selecting ref clock
    end
    // rangeA = x10 ? 5'b1 : x5 ? 5'b11110 : x2 ? 5'b10100 : x1 ? 5'b10010 : x20 ? 5'b0 : 5'b1;
    pll_rangea = 5'b00001; // 10x ref clock
    // pll_rangea = 5'b11110; // 5x ref clock
    // pll_rangea = 5'b00000; // 20x ref clock

    // JTAG simulation currently not supported here
    jtag_modesel = 1'b1;
    jtag_datain = 1'b0;

`ifndef SYNC_MUX
    async_mux = 1'b1;
`else
    async_mux = 1'b0;
`endif

    // Init JBUS model plus some ORAM stuff
    if ($test$plusargs("oram"))
    begin
`ifndef PITON_DPI
        $init_jbus_model("mem.image", 1);
`else // ifndef PITON_DPI
        init_jbus_model_call("mem.image", 1);
`endif // ifndef PITON_DPI
`ifndef METRO_CHIPSET
`ifndef __ICARUS__
        force system.chip.ctap_oram_clk_en = 1'b1;
`endif
`endif //METRO_CHIPSET
    end
    else
    begin
`ifndef PITON_DPI
        $init_jbus_model("mem.image", 0);
`else // ifndef PITON_DPI
        $display("init_jbus_model_call");
        init_jbus_model_call("mem.image", 0);
`endif // ifndef PITON_DPI
    end

    processor_offchip_noc1_valid = 0;
    processor_offchip_noc1_data  = 0;
    offchip_processor_noc1_yummy = 0;
    processor_offchip_noc2_valid = 0;
    processor_offchip_noc2_data  = 0;
    offchip_processor_noc2_yummy = 0;
    processor_offchip_noc3_valid = 0;
    processor_offchip_noc3_data  = 0;
    offchip_processor_noc3_yummy = 0;

    // Reset PLL for 100 cycles
    repeat(100)@(posedge core_ref_clk);
    pll_rst_n = 1'b1;

    // Wait for PLL lock
    wait( pll_lock == 1'b1 );

    // After 10 cycles turn on chip-level clock enable
    repeat(10)@(posedge `CHIP_INT_CLK);
    clk_en = 1'b1;

    // After 100 cycles release reset
    repeat(100)@(posedge `CHIP_INT_CLK);
    sys_rst_n = 1'b1;
    jtag_rst_l = 1'b1;

    // Wait for SRAM init
    // trin: 5000 cycles is about the lowest for 64KB L2
    // 128KB L2 requires at least 10000
    repeat(5000)@(posedge `CHIP_INT_CLK); // trin: supports at least 512KB L2 per-tile

    diag_done = 1'b1;
`ifndef METRO_CHIPSET
`ifndef PITONSYS_IOCTRL
    // Signal fake IOB to send wake up packet to first tile
    cmp_top.system.chipset.chipset_impl.ciop_fake_iob.ok_iob = 1'b1;
`endif // endif PITONSYS_IOCTRL
`endif // ifndef METRO_CHIPSET

//ok_iob = 1;

//metro code


// send data
$display("CHIPSET INITIALIZED");
@(posedge core_ref_clk);
for(int i = 0; i < 350000; i = i + 1)
begin
    #500;
// send data
    //$display("sending_chipset");
    mpi_send_data(offchip_processor_noc1_data, offchip_processor_noc1_valid, dest, rank, DATA_NOC_1);
    // send yummy
    mpi_send_yummy(processor_offchip_noc1_yummy, dest, rank, YUMMY_NOC_1);

    // send data
    mpi_send_data(offchip_processor_noc2_data, offchip_processor_noc2_valid, dest, rank, DATA_NOC_2);
    // send yummy
    mpi_send_yummy(processor_offchip_noc2_yummy, dest, rank, YUMMY_NOC_2);

    // send data
    mpi_send_data(offchip_processor_noc3_data, offchip_processor_noc3_valid, dest, rank, DATA_NOC_3);
    // send yummy
    mpi_send_yummy(processor_offchip_noc3_yummy, dest, rank, YUMMY_NOC_3);
    //$display("receiving_chipset");
    // receive data
    processor_offchip_noc1_data = mpi_receive_data(dest, valid_aux, DATA_NOC_1);
    processor_offchip_noc1_valid = valid_aux;
    // receive yummy
    offchip_processor_noc1_yummy = mpi_receive_yummy(dest, YUMMY_NOC_1);

    processor_offchip_noc2_data = mpi_receive_data(dest, valid_aux, DATA_NOC_2);
    processor_offchip_noc2_valid = valid_aux;
    // receive yummy
    offchip_processor_noc2_yummy = mpi_receive_yummy(dest, YUMMY_NOC_2);

    processor_offchip_noc3_data = mpi_receive_data(dest, valid_aux, DATA_NOC_3);
    processor_offchip_noc3_valid = valid_aux;
    // receive yummy
    offchip_processor_noc3_yummy = mpi_receive_yummy(dest, YUMMY_NOC_3);
    #500;
end
$display("Trace done: METRO_CHIPSET");
finalize();
$finish;
end
`endif

`ifdef VERILATOR
`ifndef METRO_CHIPSET
always @(posedge ok_iob) begin
    cmp_top.system.chipset.chipset_impl.ciop_fake_iob.ok_iob = 1'b1;
end
`endif // ifndef METRO_CHIPSET
`endif

////////////////////////////////////////////////////////
// SYNTHESIZABLE CHIPSET
///////////////////////////////////////////////////////

/*
integer j;
always @( posedge core_ref_clk )begin
		for(j=0;j<3;j++) begin 
			if(noc_chanel_in.valid[j] )  $display("noc%d_dat_in=%h",j,noc_chanel_in .data[j]); 
			if(noc_chanel_out.valid[j] )  $display("noc%d_dat_out=%h",j,noc_chanel_out .data[j]); 
		end
end
*/

/*
always @(posedge core_ref_clk)begin 
	if(processor_offchip_noc1_valid) $display("noc1_dat_in=%h",processor_offchip_noc1_data); 
	if(processor_offchip_noc2_valid) $display("noc2_dat_in=%h",processor_offchip_noc2_data); 
	if(processor_offchip_noc3_valid) $display("noc3_dat_in=%h",processor_offchip_noc3_data); 
	
end
*/

`ifdef PITON_PRONOC


assign smart_max = SMART_MAX;

localparam CHIP_SET_ID = T1*T2*T3+2*T1; // endp connected  of west port of router 0-0
localparam CHIP_SET_PORT = 3; //west port of first router

//off chip connection 

//NOC1
	wire [RAw-1 : 0] tile_0_0_current_r_addr1;
	wire pronoc_reset = ~sys_rst_n;
	
	
    piton_to_pronoc_wrapper #(.FLATID_WIDTH(`JTAG_FLATID_WIDTH),.NOC_NUM(1),.CHIP_SET_PORT(CHIP_SET_PORT)) pi2pr_wrapper1
	(
	.default_chipid({`NOC_CHIPID_WIDTH{1'b0}}), .default_coreid_x({`NOC_X_WIDTH{1'b0}}), .default_coreid_y({`NOC_Y_WIDTH{1'b0}}), .flat_tileid({`JTAG_FLATID_WIDTH{1'b0}}),	
	.reset(pronoc_reset),
    .clk (core_ref_clk),
	.dataIn(offchip_processor_noc1_data),
    .validIn(offchip_processor_noc1_valid),
    .yummyIn(processor_offchip_noc1_yummy),
	.chan_out(noc_chanel_out.smartflit_chanel[0]),
	.current_r_addr_i(tile_0_0_current_r_addr1)
	);	

	pronoc_to_piton_wrapper  #(.FLATID_WIDTH(`JTAG_FLATID_WIDTH),.NOC_NUM(1),.PORT_NUM(CHIP_SET_PORT)) pr2pi_wrapper1
	(
	.default_chipid({`NOC_CHIPID_WIDTH{1'b0}}), .default_coreid_x({`NOC_X_WIDTH{1'b0}}), .default_coreid_y({`NOC_Y_WIDTH{1'b0}}), .flat_tileid({`JTAG_FLATID_WIDTH{1'b0}}),	
	.reset(pronoc_reset),
    .clk (core_ref_clk),
	.dataOut(processor_offchip_noc1_data),
	.validOut(processor_offchip_noc1_valid),
	.yummyOut(offchip_processor_noc1_yummy),
	.chan_in(noc_chanel_in.smartflit_chanel[0]),
	.current_r_addr_o(tile_0_0_current_r_addr1)
	);	

//NOC2
     wire [RAw-1 : 0] tile_0_0_current_r_addr2;
    
     piton_to_pronoc_wrapper #(.FLATID_WIDTH(`JTAG_FLATID_WIDTH),.NOC_NUM(2),.CHIP_SET_PORT(CHIP_SET_PORT)) pi2pr_wrapper2
	(
	.default_chipid({`NOC_CHIPID_WIDTH{1'b0}}), .default_coreid_x({`NOC_X_WIDTH{1'b0}}), .default_coreid_y({`NOC_Y_WIDTH{1'b0}}), .flat_tileid({`JTAG_FLATID_WIDTH{1'b0}}),	
	.reset(pronoc_reset),
    .clk (core_ref_clk),
	.dataIn(offchip_processor_noc2_data),
    .validIn(offchip_processor_noc2_valid),
    .yummyIn(processor_offchip_noc2_yummy),
	.chan_out(noc_chanel_out.smartflit_chanel[1]),
	.current_r_addr_i(tile_0_0_current_r_addr2)
	);	

	pronoc_to_piton_wrapper  #(.FLATID_WIDTH(`JTAG_FLATID_WIDTH),.NOC_NUM(2),.PORT_NUM(CHIP_SET_PORT)) pr2pi_wrapper2
	(
	.default_chipid({`NOC_CHIPID_WIDTH{1'b0}}), .default_coreid_x({`NOC_X_WIDTH{1'b0}}), .default_coreid_y({`NOC_Y_WIDTH{1'b0}}), .flat_tileid({`JTAG_FLATID_WIDTH{1'b0}}),	
	.reset(pronoc_reset),
    .clk (core_ref_clk),
	.dataOut(processor_offchip_noc2_data),
	.validOut(processor_offchip_noc2_valid),
	.yummyOut(offchip_processor_noc2_yummy),
	.chan_in(noc_chanel_in.smartflit_chanel[1]),
	.current_r_addr_o(tile_0_0_current_r_addr2)
	);	


//NOC3

	wire [RAw-1 : 0] tile_0_0_current_r_addr3;

     piton_to_pronoc_wrapper #(.FLATID_WIDTH(`JTAG_FLATID_WIDTH),.NOC_NUM(3),.CHIP_SET_PORT(CHIP_SET_PORT))  pi2pr_wrapper3
	(
	.default_chipid({`NOC_CHIPID_WIDTH{1'b0}}), .default_coreid_x({`NOC_X_WIDTH{1'b0}}), .default_coreid_y({`NOC_Y_WIDTH{1'b0}}), .flat_tileid({`JTAG_FLATID_WIDTH{1'b0}}),	
	.reset(pronoc_reset),
    .clk (core_ref_clk),
	.dataIn(offchip_processor_noc3_data),
    .validIn(offchip_processor_noc3_valid),
    .yummyIn(processor_offchip_noc3_yummy),
	.chan_out(noc_chanel_out.smartflit_chanel[2]),
	.current_r_addr_i(tile_0_0_current_r_addr3)
	);	

	pronoc_to_piton_wrapper  #(.FLATID_WIDTH(`JTAG_FLATID_WIDTH),.NOC_NUM(3),.PORT_NUM(CHIP_SET_PORT)) pr2pi_wrapper3
	(
	.default_chipid({`NOC_CHIPID_WIDTH{1'b0}}), .default_coreid_x({`NOC_X_WIDTH{1'b0}}), .default_coreid_y({`NOC_Y_WIDTH{1'b0}}), .flat_tileid({`JTAG_FLATID_WIDTH{1'b0}}),	
	.reset(pronoc_reset),
    .clk (core_ref_clk),
	.dataOut(processor_offchip_noc3_data),
	.validOut(processor_offchip_noc3_valid),
	.yummyOut(offchip_processor_noc3_yummy),
	.chan_in(noc_chanel_in.smartflit_chanel[2]),
	.current_r_addr_o(tile_0_0_current_r_addr3)
	);	





`else

	assign smart_max = 0;

    assign processor_offchip_noc1_valid  =noc_chanel_in.valid [0]      ;
    assign processor_offchip_noc1_data   =noc_chanel_in.data1      ;
    assign noc_chanel_out.yummy[0]       =processor_offchip_noc1_yummy ;
                                         
    assign processor_offchip_noc2_valid  =noc_chanel_in.valid [1]      ;
    assign processor_offchip_noc2_data   =noc_chanel_in.data2      ;
    assign noc_chanel_out.yummy[1]       =processor_offchip_noc2_yummy ;
                                         
    assign processor_offchip_noc3_valid  =noc_chanel_in.valid [2]      ;
    assign processor_offchip_noc3_data   =noc_chanel_in.data3      ;
    assign noc_chanel_out.yummy[2]       =processor_offchip_noc3_yummy ;
                                         
    assign noc_chanel_out.valid[0]       =offchip_processor_noc1_valid ;
    assign noc_chanel_out.data1       =offchip_processor_noc1_data  ;
	assign offchip_processor_noc1_yummy  =noc_chanel_in.yummy [0]      ;
	                                     
	assign noc_chanel_out.valid[1]       =offchip_processor_noc2_valid ;
    assign noc_chanel_out.data2       =offchip_processor_noc2_data  ;
	assign offchip_processor_noc2_yummy  =noc_chanel_in.yummy [1]      ;
	                                     
	assign noc_chanel_out.valid[2]       =offchip_processor_noc3_valid ;
    assign noc_chanel_out.data3     =offchip_processor_noc3_data  ;
	assign offchip_processor_noc3_yummy  =noc_chanel_in.yummy [2]      ;
	
`endif
  





chipset chipset(
    .chipset_clk(core_ref_clk),

    .rst_n(sys_rst_n),

    .piton_prsnt_n(1'b0),
    .piton_ready_n(1'b0),

`ifndef PITON_BOARD
    .chipset_prsnt_n (),
`endif  // PITON_BOARD

    // Synchronous with core_ref_clk (same as io_clk in this case) and no virtual channels
    .processor_offchip_noc1_valid   (processor_offchip_noc1_valid),
    .processor_offchip_noc1_data    (processor_offchip_noc1_data),
    .processor_offchip_noc1_yummy   (processor_offchip_noc1_yummy),
    .processor_offchip_noc2_valid   (processor_offchip_noc2_valid),
    .processor_offchip_noc2_data    (processor_offchip_noc2_data),
    .processor_offchip_noc2_yummy   (processor_offchip_noc2_yummy),
    .processor_offchip_noc3_valid   (processor_offchip_noc3_valid),
    .processor_offchip_noc3_data    (processor_offchip_noc3_data),
    .processor_offchip_noc3_yummy   (processor_offchip_noc3_yummy),

    .offchip_processor_noc1_valid   (offchip_processor_noc1_valid),
    .offchip_processor_noc1_data    (offchip_processor_noc1_data),
    .offchip_processor_noc1_yummy   (offchip_processor_noc1_yummy),
    .offchip_processor_noc2_valid   (offchip_processor_noc2_valid),
    .offchip_processor_noc2_data    (offchip_processor_noc2_data),
    .offchip_processor_noc2_yummy   (offchip_processor_noc2_yummy),
    .offchip_processor_noc3_valid   (offchip_processor_noc3_valid),
    .offchip_processor_noc3_data    (offchip_processor_noc3_data),
    .offchip_processor_noc3_yummy   (offchip_processor_noc3_yummy),
    
`ifdef PITON_EXTRA_MEMS //extra mems are connected using metro_fake_mem.  
    .processor_mcx_noc2_data ( ),
    .processor_mcx_noc2_valid( ),
    .processor_mcx_noc2_yummy( ),

    .mcx_processor_noc3_data ( ),
    .mcx_processor_noc3_valid( ),
    .mcx_processor_noc3_yummy( ),
`endif
    

    // DRAM and I/O interfaces
`ifndef PITONSYS_NO_MC
`ifdef PITON_FPGA_MC_DDR3
    // FPGA DDR MC interface, currently not supported in simulation
    .init_calib_complete(),
    .ddr_addr(),
    .ddr_ba(),
    .ddr_cas_n(),
    .ddr_ck_n(),
    .ddr_ck_p(),
    .ddr_cke(),
    .ddr_ras_n(),
    .ddr_reset_n(),
    .ddr_we_n(),
    .ddr_dq(),
    .ddr_dqs_n(),
    .ddr_dqs_p(),
    .ddr_cs_n(),
    .ddr_dm(),
    .ddr_odt(),
`endif // endif PITON_FPGA_MC_DDR3
`endif // endif PITONSYS_NO_MC

`ifdef PITONSYS_IOCTRL
`ifdef PITONSYS_UART
    // UART interface for bootloading and
    // serial port interface.  Currently
    // not supported in simulation
    .uart_tx(),
    .uart_rx(),
`endif // endif PITONSYS_UART

`ifdef PITONSYS_SPI
    // SPI interface for boot device and disk.
    // Currently not supported in simulation
    .spi_data_in(),
    .spi_data_out(),
    .spi_clk_out(),
    .spi_cs_n(),
`endif // endif PITONSYS_SPI
`endif // endif PITONSYS_IOCTRL

    // Switches
`ifdef PITON_NOC_POWER_CHIPSET_TEST
    .sw({4'bz, 4'd`PITON_NOC_POWER_CHIPSET_TEST_HOP_COUNT}),
`else // ifndef PITON_NOC_POWER_CHIPSET_TEST
    .sw(),
`endif // endif PITON_NOC_POWER_CHIPSET_TEST

    // Do not provide any functionality
    .leds()

`ifdef PITON_ARIANE
    ,
    // Debug
    .ndmreset_o                     (                   ), // non-debug module reset
    .dmactive_o                     (                   ), // debug module is active
    .debug_req_o                    (                   ), // async debug request
    .unavailable_i                  ( '0                ), // communicate whether the hart is unavailable (e.g.: power down)
    // JTAG
    .tck_i                          ( '0                    ),
    .tms_i                          ( '0                    ),
    .trst_ni                        ( '0                    ),
    .td_i                           ( '0                    ),
    .td_o                           (                        ),
    .tdo_oe_o                       (                            ),
    //CLINT
    .rtc_i                          ( '0                        ), // Real-time clock in (usually 32.768 kHz)
    .timer_irq_o                    (                   ), // Timer interrupts
    .ipi_o                          (                   ), // software interrupt (a.k.a inter-process-interrupt)
    // PLIC
    .irq_o                          (                  )  // level sensitive IR lines, mip & sip (async)
`endif
`ifdef PITON_LAGARTO
    ,
    // Debug
    .ndmreset_o                     (                   ), // non-debug module reset
    .dmactive_o                     (                   ), // debug module is active
    .debug_req_o                    (                   ), // async debug request
    .unavailable_i                  ( '0                ), // communicate whether the hart is unavailable (e.g.: power down)
    // JTAG
    .tck_i                          ( '0                    ),
    .tms_i                          ( '0                    ),
    .trst_ni                        ( '0                    ),
    .td_i                           ( '0                    ),
    .td_o                           (                        ),
    .tdo_oe_o                       (                            ),
    //CLINT
    .rtc_i                          ( '0                        ), // Real-time clock in (usually 32.768 kHz)
    .timer_irq_o                    (                   ), // Timer interrupts
    .ipi_o                          (                   ), // software interrupt (a.k.a inter-process-interrupt)
    // PLIC
    .irq_o                          (                  )  // level sensitive IR lines, mip & sip (async)
`endif
);

////////////////////////////////////////////////////////
// MONITOR STUFF
////////////////////////////////////////////////////////


`ifndef DISABLE_ALL_MONITORS

    // this is the T1 sparc core monitor
    monitor   monitor(
        .clk    (`CHIP_INT_CLK),
        .cmp_gclk  (`CHIP_INT_CLK),
        .rst_l     (sys_rst_n)
        );

`ifndef MINIMAL_MONITORING

    iob_mon iob_mon(
        .clk (core_ref_clk)
    );

    integer j;

    // Tri: slam init is taken out because it's too complicated to extend to 64 cores
    // slam_init slam_init () ;

    // The only thing that we will "slam init" is the integer register file
    //  and it is randomized. For some reason if we left it as X's some tests will fail

`ifndef METRO_CHIPSET
`ifndef VERILATOR
    // T1's TSO monitor, stripped of all L2 references
    tso_mon tso_mon(`CHIP_INT_CLK, `CHIP.rst_n_inter_sync);
`endif
`endif //METRO_CHIPSET

`ifndef METRO_CHIPSET
    // L15 MONITORS
    cmp_l15_messages_mon l15_messages_mon(
        .clk (`CHIP_INT_CLK)
        );

    // DMBR MONITOR
    dmbr_mon dmbr_mon (
        .clk(`CHIP_INT_CLK)
     );

    //L2 MONITORS
    `ifdef FAKE_L2
    `else
    l2_mon l2_mon(
        .clk (`CHIP_INT_CLK)
    );
    `endif

    //only works if clk == chipset_clk
    //async_fifo_mon async_fifo_mon(
    //   .clk (core_ref_clk)
    //);

    jtag_mon jtag_mon(
        .clk (jtag_clk)
        );

    iob_mon iob_mon(
        .clk (chipset_clk)
    );
    // sas, more debug info
`endif // ifndef METRO_CHIPSET

    // turn on sas interface after a delay
//    reg   need_sas_sparc_intf_update;
//    initial begin
//        need_sas_sparc_intf_update  = 0;
//        #12500;
//        need_sas_sparc_intf_update  = 1;
//    end // initial begin

`ifdef PITON_OST1
    sas_intf  sas_intf(/*AUTOINST*/
        // Inputs
        .clk       (`CHIP_INT_CLK),      // Templated
        .rst_l     (`CHIP.rst_n_inter_sync));       // Templated
`endif

`ifdef PITON_OST1
    // create sas tasks
    sas_tasks sas_tasks(/*AUTOINST*/
        // Inputs
        .clk      (`CHIP_INT_CLK),      // Templated
        .rst_l        (`CHIP.rst_n_inter_sync));       // Templated
`endif

`ifdef PITON_OST1
    // sparc pipe flow monitor
    sparc_pipe_flow sparc_pipe_flow(/*AUTOINST*/
        // Inputs
        .clk  (`CHIP_INT_CLK));         // Templated
`endif

`ifndef METRO_CHIPSET
    manycore_network_mon network_mon (`CHIP_INT_CLK);
`endif // ifndef METRO_CHIPSET

`endif // MINIMAL_MONITORING
`endif // DISABLE_ALL_MONITORS
    // Alexey
    // UART monitor
    /*reg      prev_tx_state;
    always @(posedge core_ref_clk)
        prev_tx_state <= tx;

    always @(posedge core_ref_clk)
        if (prev_tx_state != tx) begin
            $display("UART: TX changed to %d at", tx, $time);
        end*/



`ifdef VERILATOR
`ifdef METRO_CHIPSET


`define MY_CHIPSET  `TOP_MOD_INST.chipset_impl 
 test_end_checker test_end_checker(
            .clk                    (`MY_CHIPSET.chipset_clk),
            .rst_n                  (`MY_CHIPSET.chipset_rst_n),

            .src_checker_noc2_val   (`MY_CHIPSET.chip_filter_noc2_valid),
            .src_checker_noc2_data  (`MY_CHIPSET.chip_filter_noc2_data),
            .src_checker_noc2_rdy   (`MY_CHIPSET.filter_chip_noc2_ready),

            .uart_boot_en           (test_ena),
            .test_good_end          (good_end),
            .test_bad_end           (bad_end)
        );
 
`endif // METRO_CHIPSET

    assign flit_o_cnts=`MY_CHIPSET.fake_mem_ctrl.flit_o_cnts;
    assign flit_i_cnts=`MY_CHIPSET.fake_mem_ctrl.flit_i_cnts;

`endif // VERILATOR


endmodule // cmp_top

`endif
